module start_sprite_control(
	input clk,
	input draw,
    input clear,
    input shift_h,
    input shift_v,
    input load,
    input [6:0] shift_amount,
    input [7:0] load_x,
    input [6:0] load_y,
    output reg complete,
    output reg [7:0] x_out,
    output reg [6:0] y_out,
    output reg [11:0] colour_out,
    output reg [7:0] posx,
    output reg [6:0] posy
    );

    reg [7:0] x_pos;
    reg [6:0] y_pos;
    reg [11:0] sprite [0:511]; 
    reg [8:0] pointer;

    initial begin
        x_pos = 8'd49;
        y_pos = 7'd48;
        pointer = 1'b1;

        sprite[0] = 12'b000000000000;
        sprite[1] = 12'b000000000000;
        sprite[2] = 12'b000000000000;
        sprite[3] = 12'b000000000000;
        sprite[4] = 12'b000000000000;
        sprite[5] = 12'b000000000000;
        sprite[6] = 12'b000000000000;
        sprite[7] = 12'b000000000000;
        sprite[8] = 12'b000000000000;
        sprite[9] = 12'b000000000000;
        sprite[10] = 12'b000000000000;
        sprite[11] = 12'b000000000000;
        sprite[12] = 12'b000000000000;
        sprite[13] = 12'b000000000000;
        sprite[14] = 12'b000000000000;
        sprite[15] = 12'b000000000000;
        sprite[16] = 12'b000000000000;
        sprite[17] = 12'b000000000000;
        sprite[18] = 12'b000000000000;
        sprite[19] = 12'b000000000000;
        sprite[20] = 12'b000000000000;
        sprite[21] = 12'b000000000000;
        sprite[22] = 12'b000000000000;
        sprite[23] = 12'b000000000000;
        sprite[24] = 12'b000000000000;
        sprite[25] = 12'b000000000000;
        sprite[26] = 12'b000000000000;
        sprite[27] = 12'b000000000000;
        sprite[28] = 12'b000000000000;
        sprite[29] = 12'b000000000000;
        sprite[30] = 12'b000000000000;
        sprite[31] = 12'b000000000000;
        sprite[32] = 12'b000000000000;
        sprite[33] = 12'b000000000000;
        sprite[34] = 12'b000000000000;
        sprite[35] = 12'b000000000000;
        sprite[36] = 12'b000000000000;
        sprite[37] = 12'b000000000000;
        sprite[38] = 12'b000000000000;
        sprite[39] = 12'b000000000000;
        sprite[40] = 12'b000000000000;
        sprite[41] = 12'b000000000000;
        sprite[42] = 12'b000000000000;
        sprite[43] = 12'b000000000000;
        sprite[44] = 12'b000000000000;
        sprite[45] = 12'b000000000000;
        sprite[46] = 12'b000000000000;
        sprite[47] = 12'b000000000000;
        sprite[48] = 12'b000000000000;
        sprite[49] = 12'b000000000000;
        sprite[50] = 12'b000000000000;
        sprite[51] = 12'b000000000000;
        sprite[52] = 12'b000000000000;
        sprite[53] = 12'b000000000000;
        sprite[54] = 12'b000000000000;
        sprite[55] = 12'b000000000000;
        sprite[56] = 12'b000000000000;
        sprite[57] = 12'b000000000000;
        sprite[58] = 12'b000000000000;
        sprite[59] = 12'b000000000000;
        sprite[60] = 12'b000000000000;
        sprite[61] = 12'b000000000000;
        sprite[62] = 12'b000000000000;
        sprite[63] = 12'b000000000000;
        sprite[64] = 12'b000000001111;
        sprite[65] = 12'b111111111111;
        sprite[66] = 12'b111111110000;
        sprite[67] = 12'b000000000000;
        sprite[68] = 12'b000000001111;
        sprite[69] = 12'b111111110000;
        sprite[70] = 12'b000000000000;
        sprite[71] = 12'b000000000000;
        sprite[72] = 12'b000000000000;
        sprite[73] = 12'b000000000000;
        sprite[74] = 12'b000000000000;
        sprite[75] = 12'b000000000000;
        sprite[76] = 12'b000000000000;
        sprite[77] = 12'b000000000000;
        sprite[78] = 12'b000000000000;
        sprite[79] = 12'b000000000000;
        sprite[80] = 12'b000000000000;
        sprite[81] = 12'b000000000000;
        sprite[82] = 12'b000000000000;
        sprite[83] = 12'b000000000000;
        sprite[84] = 12'b000000000000;
        sprite[85] = 12'b000000000000;
        sprite[86] = 12'b000000000000;
        sprite[87] = 12'b000000000000;
        sprite[88] = 12'b000000000000;
        sprite[89] = 12'b000000000000;
        sprite[90] = 12'b000000000000;
        sprite[91] = 12'b000000000000;
        sprite[92] = 12'b000000001111;
        sprite[93] = 12'b111111111111;
        sprite[94] = 12'b111111110000;
        sprite[95] = 12'b000000000000;
        sprite[96] = 12'b000000000000;
        sprite[97] = 12'b000000000000;
        sprite[98] = 12'b000000000000;
        sprite[99] = 12'b000000000000;
        sprite[100] = 12'b000000000000;
        sprite[101] = 12'b000000000000;
        sprite[102] = 12'b000000000000;
        sprite[103] = 12'b000000000000;
        sprite[104] = 12'b000000000000;
        sprite[105] = 12'b000000000000;
        sprite[106] = 12'b000000000000;
        sprite[107] = 12'b000000000000;
        sprite[108] = 12'b000000000000;
        sprite[109] = 12'b000000000000;
        sprite[110] = 12'b000000000000;
        sprite[111] = 12'b000000000000;
        sprite[112] = 12'b000000000000;
        sprite[113] = 12'b000000000000;
        sprite[114] = 12'b000000000000;
        sprite[115] = 12'b000000000000;
        sprite[116] = 12'b000000000000;
        sprite[117] = 12'b000000000000;
        sprite[118] = 12'b000000000000;
        sprite[119] = 12'b000000000000;
        sprite[120] = 12'b000000000000;
        sprite[121] = 12'b000000000000;
        sprite[122] = 12'b000000000000;
        sprite[123] = 12'b000000000000;
        sprite[124] = 12'b000000000000;
        sprite[125] = 12'b000000000000;
        sprite[126] = 12'b000000000000;
        sprite[127] = 12'b000000000000;
        sprite[128] = 12'b000000001111;
        sprite[129] = 12'b111111110000;
        sprite[130] = 12'b000000001111;
        sprite[131] = 12'b111111110000;
        sprite[132] = 12'b000000001111;
        sprite[133] = 12'b111111110000;
        sprite[134] = 12'b000000000000;
        sprite[135] = 12'b000000000000;
        sprite[136] = 12'b000000000000;
        sprite[137] = 12'b000000000000;
        sprite[138] = 12'b000000000000;
        sprite[139] = 12'b000000000000;
        sprite[140] = 12'b000000000000;
        sprite[141] = 12'b000000000000;
        sprite[142] = 12'b000000000000;
        sprite[143] = 12'b000000000000;
        sprite[144] = 12'b000000000000;
        sprite[145] = 12'b000000000000;
        sprite[146] = 12'b000000001111;
        sprite[147] = 12'b111111110000;
        sprite[148] = 12'b000000000000;
        sprite[149] = 12'b000000000000;
        sprite[150] = 12'b000000000000;
        sprite[151] = 12'b000000000000;
        sprite[152] = 12'b000000000000;
        sprite[153] = 12'b000000000000;
        sprite[154] = 12'b000000000000;
        sprite[155] = 12'b000000001111;
        sprite[156] = 12'b111111110000;
        sprite[157] = 12'b000000000000;
        sprite[158] = 12'b000000000000;
        sprite[159] = 12'b000000001111;
        sprite[160] = 12'b111111110000;
        sprite[161] = 12'b000000000000;
        sprite[162] = 12'b000000000000;
        sprite[163] = 12'b000000000000;
        sprite[164] = 12'b000000000000;
        sprite[165] = 12'b000000000000;
        sprite[166] = 12'b000000000000;
        sprite[167] = 12'b000000000000;
        sprite[168] = 12'b000000000000;
        sprite[169] = 12'b000000000000;
        sprite[170] = 12'b000000000000;
        sprite[171] = 12'b000000001111;
        sprite[172] = 12'b111111110000;
        sprite[173] = 12'b000000000000;
        sprite[174] = 12'b000000000000;
        sprite[175] = 12'b000000000000;
        sprite[176] = 12'b000000000000;
        sprite[177] = 12'b000000000000;
        sprite[178] = 12'b000000000000;
        sprite[179] = 12'b000000000000;
        sprite[180] = 12'b000000000000;
        sprite[181] = 12'b000000000000;
        sprite[182] = 12'b000000000000;
        sprite[183] = 12'b000000000000;
        sprite[184] = 12'b000000000000;
        sprite[185] = 12'b000000000000;
        sprite[186] = 12'b000000000000;
        sprite[187] = 12'b000000000000;
        sprite[188] = 12'b000000000000;
        sprite[189] = 12'b000000000000;
        sprite[190] = 12'b000000000000;
        sprite[191] = 12'b000000000000;
        sprite[192] = 12'b000000001111;
        sprite[193] = 12'b111111110000;
        sprite[194] = 12'b000000001111;
        sprite[195] = 12'b111111110000;
        sprite[196] = 12'b000000001111;
        sprite[197] = 12'b111111110000;
        sprite[198] = 12'b000000000000;
        sprite[199] = 12'b000000000000;
        sprite[200] = 12'b000000000000;
        sprite[201] = 12'b000000000000;
        sprite[202] = 12'b000000000000;
        sprite[203] = 12'b000000000000;
        sprite[204] = 12'b000000000000;
        sprite[205] = 12'b000000000000;
        sprite[206] = 12'b000000000000;
        sprite[207] = 12'b000000000000;
        sprite[208] = 12'b000000000000;
        sprite[209] = 12'b000000000000;
        sprite[210] = 12'b000000001111;
        sprite[211] = 12'b111111110000;
        sprite[212] = 12'b000000000000;
        sprite[213] = 12'b000000000000;
        sprite[214] = 12'b000000000000;
        sprite[215] = 12'b000000000000;
        sprite[216] = 12'b000000000000;
        sprite[217] = 12'b000000000000;
        sprite[218] = 12'b000000000000;
        sprite[219] = 12'b000000001111;
        sprite[220] = 12'b111111110000;
        sprite[221] = 12'b000000000000;
        sprite[222] = 12'b000000000000;
        sprite[223] = 12'b000000001111;
        sprite[224] = 12'b111111110000;
        sprite[225] = 12'b000000000000;
        sprite[226] = 12'b000000000000;
        sprite[227] = 12'b000000000000;
        sprite[228] = 12'b000000000000;
        sprite[229] = 12'b000000000000;
        sprite[230] = 12'b000000000000;
        sprite[231] = 12'b000000000000;
        sprite[232] = 12'b000000000000;
        sprite[233] = 12'b000000000000;
        sprite[234] = 12'b000000000000;
        sprite[235] = 12'b000000001111;
        sprite[236] = 12'b111111110000;
        sprite[237] = 12'b000000000000;
        sprite[238] = 12'b000000000000;
        sprite[239] = 12'b000000000000;
        sprite[240] = 12'b000000000000;
        sprite[241] = 12'b000000000000;
        sprite[242] = 12'b000000000000;
        sprite[243] = 12'b000000000000;
        sprite[244] = 12'b000000000000;
        sprite[245] = 12'b000000000000;
        sprite[246] = 12'b000000000000;
        sprite[247] = 12'b000000000000;
        sprite[248] = 12'b000000000000;
        sprite[249] = 12'b000000000000;
        sprite[250] = 12'b000000000000;
        sprite[251] = 12'b000000000000;
        sprite[252] = 12'b000000000000;
        sprite[253] = 12'b000000000000;
        sprite[254] = 12'b000000000000;
        sprite[255] = 12'b000000000000;
        sprite[256] = 12'b000000001111;
        sprite[257] = 12'b111111111111;
        sprite[258] = 12'b111111110000;
        sprite[259] = 12'b000000000000;
        sprite[260] = 12'b000000001111;
        sprite[261] = 12'b111111110000;
        sprite[262] = 12'b000000001111;
        sprite[263] = 12'b111111111111;
        sprite[264] = 12'b111111111111;
        sprite[265] = 12'b111111110000;
        sprite[266] = 12'b000000001111;
        sprite[267] = 12'b111111110000;
        sprite[268] = 12'b000000000000;
        sprite[269] = 12'b000000000000;
        sprite[270] = 12'b000000001111;
        sprite[271] = 12'b111111110000;
        sprite[272] = 12'b000000000000;
        sprite[273] = 12'b000000000000;
        sprite[274] = 12'b000000001111;
        sprite[275] = 12'b111111111111;
        sprite[276] = 12'b111111110000;
        sprite[277] = 12'b000000001111;
        sprite[278] = 12'b111111111111;
        sprite[279] = 12'b111111111111;
        sprite[280] = 12'b111111110000;
        sprite[281] = 12'b000000000000;
        sprite[282] = 12'b000000000000;
        sprite[283] = 12'b000000000000;
        sprite[284] = 12'b000000001111;
        sprite[285] = 12'b111111111111;
        sprite[286] = 12'b111111110000;
        sprite[287] = 12'b000000001111;
        sprite[288] = 12'b111111111111;
        sprite[289] = 12'b111111110000;
        sprite[290] = 12'b000000001111;
        sprite[291] = 12'b111111111111;
        sprite[292] = 12'b111111111111;
        sprite[293] = 12'b111111110000;
        sprite[294] = 12'b000000000000;
        sprite[295] = 12'b000000000000;
        sprite[296] = 12'b000000001111;
        sprite[297] = 12'b111111111111;
        sprite[298] = 12'b111111110000;
        sprite[299] = 12'b000000001111;
        sprite[300] = 12'b111111111111;
        sprite[301] = 12'b111111110000;
        sprite[302] = 12'b000000000000;
        sprite[303] = 12'b000000000000;
        sprite[304] = 12'b000000000000;
        sprite[305] = 12'b000000000000;
        sprite[306] = 12'b000000000000;
        sprite[307] = 12'b000000000000;
        sprite[308] = 12'b000000000000;
        sprite[309] = 12'b000000000000;
        sprite[310] = 12'b000000000000;
        sprite[311] = 12'b000000000000;
        sprite[312] = 12'b000000000000;
        sprite[313] = 12'b000000000000;
        sprite[314] = 12'b000000000000;
        sprite[315] = 12'b000000000000;
        sprite[316] = 12'b000000000000;
        sprite[317] = 12'b000000000000;
        sprite[318] = 12'b000000000000;
        sprite[319] = 12'b000000000000;
        sprite[320] = 12'b000000001111;
        sprite[321] = 12'b111111110000;
        sprite[322] = 12'b000000001111;
        sprite[323] = 12'b111111110000;
        sprite[324] = 12'b000000001111;
        sprite[325] = 12'b111111110000;
        sprite[326] = 12'b000000001111;
        sprite[327] = 12'b111111110000;
        sprite[328] = 12'b000000001111;
        sprite[329] = 12'b111111110000;
        sprite[330] = 12'b000000001111;
        sprite[331] = 12'b111111110000;
        sprite[332] = 12'b000000001111;
        sprite[333] = 12'b111111110000;
        sprite[334] = 12'b000000001111;
        sprite[335] = 12'b111111110000;
        sprite[336] = 12'b000000000000;
        sprite[337] = 12'b000000000000;
        sprite[338] = 12'b000000001111;
        sprite[339] = 12'b111111110000;
        sprite[340] = 12'b000000000000;
        sprite[341] = 12'b000000001111;
        sprite[342] = 12'b111111110000;
        sprite[343] = 12'b000000001111;
        sprite[344] = 12'b111111110000;
        sprite[345] = 12'b000000000000;
        sprite[346] = 12'b000000000000;
        sprite[347] = 12'b000000000000;
        sprite[348] = 12'b000000000000;
        sprite[349] = 12'b000000001111;
        sprite[350] = 12'b111111110000;
        sprite[351] = 12'b000000001111;
        sprite[352] = 12'b111111110000;
        sprite[353] = 12'b000000000000;
        sprite[354] = 12'b000000001111;
        sprite[355] = 12'b111111110000;
        sprite[356] = 12'b000000001111;
        sprite[357] = 12'b111111110000;
        sprite[358] = 12'b000000000000;
        sprite[359] = 12'b000000001111;
        sprite[360] = 12'b111111110000;
        sprite[361] = 12'b000000000000;
        sprite[362] = 12'b000000000000;
        sprite[363] = 12'b000000001111;
        sprite[364] = 12'b111111110000;
        sprite[365] = 12'b000000000000;
        sprite[366] = 12'b000000000000;
        sprite[367] = 12'b000000000000;
        sprite[368] = 12'b000000000000;
        sprite[369] = 12'b000000000000;
        sprite[370] = 12'b000000000000;
        sprite[371] = 12'b000000000000;
        sprite[372] = 12'b000000000000;
        sprite[373] = 12'b000000000000;
        sprite[374] = 12'b000000000000;
        sprite[375] = 12'b000000000000;
        sprite[376] = 12'b000000000000;
        sprite[377] = 12'b000000000000;
        sprite[378] = 12'b000000000000;
        sprite[379] = 12'b000000000000;
        sprite[380] = 12'b000000000000;
        sprite[381] = 12'b000000000000;
        sprite[382] = 12'b000000000000;
        sprite[383] = 12'b000000000000;
        sprite[384] = 12'b000000001111;
        sprite[385] = 12'b111111111111;
        sprite[386] = 12'b111111110000;
        sprite[387] = 12'b000000000000;
        sprite[388] = 12'b000000001111;
        sprite[389] = 12'b111111110000;
        sprite[390] = 12'b000000001111;
        sprite[391] = 12'b111111111111;
        sprite[392] = 12'b111111111111;
        sprite[393] = 12'b111111110000;
        sprite[394] = 12'b000000000000;
        sprite[395] = 12'b000000001111;
        sprite[396] = 12'b111111110000;
        sprite[397] = 12'b000000001111;
        sprite[398] = 12'b111111110000;
        sprite[399] = 12'b000000000000;
        sprite[400] = 12'b000000000000;
        sprite[401] = 12'b000000000000;
        sprite[402] = 12'b000000001111;
        sprite[403] = 12'b111111111111;
        sprite[404] = 12'b111111110000;
        sprite[405] = 12'b000000001111;
        sprite[406] = 12'b111111111111;
        sprite[407] = 12'b111111111111;
        sprite[408] = 12'b111111110000;
        sprite[409] = 12'b000000000000;
        sprite[410] = 12'b000000000000;
        sprite[411] = 12'b000000001111;
        sprite[412] = 12'b111111111111;
        sprite[413] = 12'b111111110000;
        sprite[414] = 12'b000000000000;
        sprite[415] = 12'b000000001111;
        sprite[416] = 12'b111111111111;
        sprite[417] = 12'b111111110000;
        sprite[418] = 12'b000000001111;
        sprite[419] = 12'b111111111111;
        sprite[420] = 12'b111111110000;
        sprite[421] = 12'b000000001111;
        sprite[422] = 12'b111111110000;
        sprite[423] = 12'b000000001111;
        sprite[424] = 12'b111111110000;
        sprite[425] = 12'b000000000000;
        sprite[426] = 12'b000000000000;
        sprite[427] = 12'b000000001111;
        sprite[428] = 12'b111111111111;
        sprite[429] = 12'b111111110000;
        sprite[430] = 12'b000000000000;
        sprite[431] = 12'b000000000000;
        sprite[432] = 12'b000000000000;
        sprite[433] = 12'b000000000000;
        sprite[434] = 12'b000000000000;
        sprite[435] = 12'b000000000000;
        sprite[436] = 12'b000000000000;
        sprite[437] = 12'b000000000000;
        sprite[438] = 12'b000000000000;
        sprite[439] = 12'b000000000000;
        sprite[440] = 12'b000000000000;
        sprite[441] = 12'b000000000000;
        sprite[442] = 12'b000000000000;
        sprite[443] = 12'b000000000000;
        sprite[444] = 12'b000000000000;
        sprite[445] = 12'b000000000000;
        sprite[446] = 12'b000000000000;
        sprite[447] = 12'b000000000000;
        sprite[448] = 12'b000000000000;
        sprite[449] = 12'b000000000000;
        sprite[450] = 12'b000000000000;
        sprite[451] = 12'b000000000000;
        sprite[452] = 12'b000000000000;
        sprite[453] = 12'b000000000000;
        sprite[454] = 12'b000000000000;
        sprite[455] = 12'b000000000000;
        sprite[456] = 12'b000000000000;
        sprite[457] = 12'b000000000000;
        sprite[458] = 12'b000000000000;
        sprite[459] = 12'b000000000000;
        sprite[460] = 12'b000000000000;
        sprite[461] = 12'b000000000000;
        sprite[462] = 12'b000000000000;
        sprite[463] = 12'b000000000000;
        sprite[464] = 12'b000000000000;
        sprite[465] = 12'b000000000000;
        sprite[466] = 12'b000000000000;
        sprite[467] = 12'b000000000000;
        sprite[468] = 12'b000000000000;
        sprite[469] = 12'b000000000000;
        sprite[470] = 12'b000000000000;
        sprite[471] = 12'b000000000000;
        sprite[472] = 12'b000000000000;
        sprite[473] = 12'b000000000000;
        sprite[474] = 12'b000000000000;
        sprite[475] = 12'b000000000000;
        sprite[476] = 12'b000000000000;
        sprite[477] = 12'b000000000000;
        sprite[478] = 12'b000000000000;
        sprite[479] = 12'b000000000000;
        sprite[480] = 12'b000000000000;
        sprite[481] = 12'b000000000000;
        sprite[482] = 12'b000000000000;
        sprite[483] = 12'b000000000000;
        sprite[484] = 12'b000000000000;
        sprite[485] = 12'b000000000000;
        sprite[486] = 12'b000000000000;
        sprite[487] = 12'b000000000000;
        sprite[488] = 12'b000000000000;
        sprite[489] = 12'b000000000000;
        sprite[490] = 12'b000000000000;
        sprite[491] = 12'b000000000000;
        sprite[492] = 12'b000000000000;
        sprite[493] = 12'b000000000000;
        sprite[494] = 12'b000000000000;
        sprite[495] = 12'b000000000000;
        sprite[496] = 12'b000000000000;
        sprite[497] = 12'b000000000000;
        sprite[498] = 12'b000000000000;
        sprite[499] = 12'b000000000000;
        sprite[500] = 12'b000000000000;
        sprite[501] = 12'b000000000000;
        sprite[502] = 12'b000000000000;
        sprite[503] = 12'b000000000000;
        sprite[504] = 12'b000000000000;
        sprite[505] = 12'b000000000000;
        sprite[506] = 12'b000000000000;
        sprite[507] = 12'b000000000000;
        sprite[508] = 12'b000000000000;
        sprite[509] = 12'b000000000000;
        sprite[510] = 12'b000000000000;
        sprite[511] = 12'b000000000000;
    end

    always@(negedge clk) begin
		  if (draw) begin
			  if (clear) 
					begin
						 x_out = x_pos + pointer[5:0];
						 y_out = y_pos + pointer[8:6];
						 colour_out = 1'b0;
						 pointer = pointer + 1'b1;
					end
			  else if (shift_h)
					begin
						 // x_out = x_pos + shift_amount + pointer[5:0];
						 x_out = x_pos + pointer[5:0];
						 y_out = y_pos + pointer[8:6];
						 colour_out = sprite[pointer];
						 pointer = pointer + 1'b1;
//						 if (pointer == 1'b0)
//							  x_pos = x_pos + shift_amount;
					end
//			  else if (shift_v)
//					begin
//						 x_out = x_pos + pointer[5:0];
//						 y_out = y_pos + shift_amount + pointer[8:6];
//						 colour_out = sprite[pointer];
//						 pointer = pointer + 1'b1;
//						 if (pointer == 1'b0)
//							  y_pos = y_pos + shift_amount;
//					end
//            else if (load)
//                begin
//                    x_pos = load_x;
//                    y_pos = load_y;
//                end
		end
    end

    always @(*)begin
		if(pointer == 1'b0)
		begin
			complete = 1'b1;
			posy <= y_pos;
			posx <= x_pos;
		end
		else
			complete = 1'b0;
	end
endmodule